.subckt cpw a b p len=220u width=4.4u space=4.4u scale=0.90909090909091
*
.param
*
+ l = '(len*scale)'
+ w = '(width*scale)*1e6'
+ s = '(space*scale)*1e6'
*
*
+ R0_unit = '((5.401614077061407e3)+(-1.169578893808857e3)*w+(-1.514201973460804e2)*s+(1.320756713699097e2)*(w**2)+(-1.380780197344119e1)*w*s+(2.869594793526634e1)*(s**2)+(-5.197930007226441)*(w**3)+(4.411520322137612e-1)*(w**2)*s+(6.159679369564878e-1)*w*(s**2)+(-1.597137968961264)*(s**3))'
+ R1_unit = '((3.109803805636977e2)+(-2.133728103009985e1)*w+(-4.947659839352988e1)*s+(2.317684449970950e1)*(w**2)+(-3.262165464371888e1)*w*s+(2.251320853316543e1)*(s**2)+(-1.526242680760257)*(w**3)+(1.065331535849124)*(w**2)*s+(1.072233639045007)*w*(s**2)+(-1.407697001476457)*(s**3))'
+ R2_unit = '((7.838554776552836e3)+(8.003075897531999e2)*w+(-2.104465732866399e3)*s+(-1.507068951177143e2)*(w**2)+(6.128293705828987e1)*w*s+(2.654002598018084e2)*(s**2)+(5.050859953171345)*(w**3)+(3.937300359713792)*(w**2)*s+(-8.828719921808693)*w*(s**2)+(-9.112573329000233)*(s**3))'
+ R3_unit = '((3.220338406646986e3)+(-2.489958997643127e3)*w+(4.875972775109543e3)*s+(1.398313480753162e2)*(w**2)+(2.526769350075681e2)*w*s+(-8.547690905398572e2)*(s**2)+(1.235736934955830)*(w**3)+(-1.241623247096959e1)*(w**2)*s+(-5.259446001007047)*w*(s**2)+(4.229939671650986e1)*(s**3))'
+ L0_unit = '((1.685484858516990e-7)+(-2.249123501494398e-8)*w+(5.934432147440323e-8)*s+(3.251379216964253e-9)*(w**2)+(-4.095410448197849e-9)*w*s+(-1.296219748327626e-9)*(s**2)+(-1.555462582632252e-10)*(w**3)+(1.352600972914807e-10)*(w**2)*s+(1.152935734969073e-10)*w*(s**2)+(-3.891285683439306e-11)*(s**3))'
+ L1_unit = '((4.949406477131133e-8)+(-3.395933748081339e-9)*w+(-7.874445201702794e-9)*s+(3.688709367400977e-9)*(w**2)+(-5.191897588384542e-9)*w*s+(3.583088422911913e-9)*(s**2)+(-2.429090670008207e-10)*(w**3)+(1.695527799620688e-10)*(w**2)*s+(1.706512838034240e-10)*w*(s**2)+(-2.240419361606170e-10)*(s**3))'
+ L2_unit = '((5.100388690735639e-8)+(-8.477728692172104e-10)*w+(-4.381830106951298e-9)*s+(-6.837810032587059e-10)*(w**2)+(1.690700339947600e-9)*w*s+(-1.692800554800766e-10)*(s**2)+(5.222326237810560e-11)*(w**3)+(-6.312708500390784e-11)*(w**2)*s+(-5.886496808760335e-11)*w*(s**2)+(3.077424835881944e-11)*(s**3))'
+ L3_unit = '((5.125327758465446e-9)+(-3.962892825710448e-9)*w+(7.760351695401912e-9)*s+(2.225485024538999e-10)*(w**2)+(4.021478321176401e-10)*w*s+(-1.360407259615822e-9)*(s**2)+(1.966736415594459e-12)*(w**3)+(-1.976104772332907e-11)*(w**2)*s+(-8.370668289851722e-12)*w*(s**2)+(6.732158077237638e-11)*(s**3))'
+ G0_unit = '((-5.564365322650253e-2)+(1.693710631950140e-2)*w+(1.172803173649778e-2)*s+(-1.786992046156378e-3)*(w**2)+(-1.647724334506544e-3)*w*s+(-8.829040066258833e-4)*(s**2)+(7.745084450107837e-5)*(w**3)+(7.499115309252783e-5)*(w**2)*s+(6.967431040567679e-5)*w*(s**2)+(2.400150856927265e-5)*(s**3))'
+ G1_unit = '((8.973701959700016e-2)+(-2.896735110684835e-2)*w+(-2.230938096092836e-2)*s+(2.925618632752435e-3)*(w**2)+(4.253215862929393e-3)*w*s+(2.024138928091936e-3)*(s**2)+(-1.093240263227041e-4)*(w**3)+(-1.382091102680441e-4)*(w**2)*s+(-1.628911975255663e-4)*w*(s**2)+(-5.609493494529538e-5)*(s**3))'
+ G2_unit = '((-1.021426894417850)+(1.010669419336415e-1)*w+(2.585712658212557e-1)*s+(-4.490868214944547e-3)*(w**2)+(1.952999739605092e-2)*w*s+(-2.422759952917492e-2)*(s**2)+(4.341981885288029e-4)*(w**3)+(-9.093745277283890e-4)*(w**2)*s+(-3.785289550046849e-4)*w*(s**2)+(1.002705667192365e-3)*(s**3))'
+ G3_unit = '((2.544068912925331)+(-1.329244621135182e-1)*w+(-8.063053013408309e-1)*s+(2.073833313033228e-2)*(w**2)+(-6.217774535397997e-3)*w*s+(1.062121477597713e-1)*(s**2)+(-9.354851741958824e-4)*(w**3)+(7.600451481945094e-4)*(w**2)*s+(-1.469604562330072e-4)*w*(s**2)+(-4.599480542243937e-3)*(s**3))'
+ C0_unit = '((3.083615389585745e-10)+(1.284756028574325e-11)*w+(-6.896593157690734e-11)*s+(-5.025935494630162e-13)*(w**2)+(-9.976350598510736e-13)*w*s+(7.662011432148645e-12)*(s**2)+(1.273669644571410e-14)*(w**3)+(1.945878824590009e-14)*(w**2)*s+(3.727114000946531e-14)*w*(s**2)+(-3.031328557138464e-13)*(s**3))'
+ C1_unit = '((1.428209024719684e-11)+(-4.610297116933401e-12)*w+(-3.550648257251963e-12)*s+(4.656266670043025e-13)*(w**2)+(6.769203286220741e-13)*w*s+(3.221517159105616e-13)*(s**2)+(-1.739945918796684e-14)*(w**3)+(-2.199666307949205e-14)*(w**2)*s+(-2.592493927235217e-14)*w*(s**2)+(-8.927786178962044e-15)*(s**3))'
+ C2_unit = '((-1.509020342826772e-11)+(2.711214390797377e-12)*w+(2.873172936234656e-12)*s+(-2.708056993196995e-13)*(w**2)+(2.478040765466568e-13)*w*s+(-2.092989056952832e-13)*(s**2)+(1.702142825426101e-14)*(w**3)+(-4.213984931156892e-15)*(w**2)*s+(-4.568413842642727e-15)*w*(s**2)+(8.631113579411743e-15)*(s**3))'
+ C3_unit = '((4.049011430584910e-12)+(-2.115558520319776e-13)*w+(-1.283274743495934e-12)*s+(3.300608229178798e-14)*(w**2)+(-9.895895523395049e-15)*w*s+(1.690418833237438e-13)*(s**2)+(-1.488870896624573e-15)*(w**3)+(1.209649423081684e-15)*(w**2)*s+(-2.338948304852326e-16)*w*(s**2)+(-7.320300639531133e-15)*(s**3))'
*
+ R0  = 'l*R0_unit/10'
+ R1  = 'l*R1_unit/10'
+ R2  = 'l*R2_unit/10'
+ R3  = 'l*R3_unit/10'
+ L0  = 'l*L0_unit/10'
+ L1  = 'l*L1_unit/10'
+ L2  = 'l*L2_unit/10'
+ L3  = 'l*L3_unit/10'
+ RG0 = '10/(l*G0_unit)'
+ RG1 = '10/(l*G1_unit)'
+ RG2 = '10/(l*G2_unit)'
+ RG3 = '10/(l*G3_unit)'
+ C0  = 'l*C0_unit/10'
+ C1  = 'l*C1_unit/10'
+ C2  = 'l*C2_unit/10'
+ C3  = 'l*C3_unit/10'
*
*
*
*******************************************************
******                  Netlist                  ******
*******************************************************
RG010      		a          		p          		'2*RG0'
C010       		a          		p          		'0.5*C0'
RG011      		a          		np011      		'2*RG1'
C011       		np011      		p          		'0.5*C1'
RG012      		a          		np012      		'2*RG2'
C012       		np012      		p          		'0.5*C2'
RG013      		a          		np013      		'2*RG3'
C013       		np013      		p          		'0.5*C3'
R010       		a          		ns011      		'R0'
L010       		ns011      		ns012      		'L0'
R011       		ns012      		ns013      		'R1'
L011       		ns012      		ns013      		'L1'
R012       		ns013      		ns014      		'R2'
L012       		ns013      		ns014      		'L2'
R013       		ns014      		ns015      		'R3'
L013       		ns014      		ns015      		'L3'
RG020      		ns015      		p          		'RG0'
C020       		ns015      		p          		'C0'
RG021      		ns015      		np021      		'RG1'
C021       		np021      		p          		'C1'
RG022      		ns015      		np022      		'RG2'
C022       		np022      		p          		'C2'
RG023      		ns015      		np023      		'RG3'
C023       		np023      		p          		'C3'
R020       		ns015      		ns021      		'R0'
L020       		ns021      		ns022      		'L0'
R021       		ns022      		ns023      		'R1'
L021       		ns022      		ns023      		'L1'
R022       		ns023      		ns024      		'R2'
L022       		ns023      		ns024      		'L2'
R023       		ns024      		ns025      		'R3'
L023       		ns024      		ns025      		'L3'
RG030      		ns025      		p          		'RG0'
C030       		ns025      		p          		'C0'
RG031      		ns025      		np031      		'RG1'
C031       		np031      		p          		'C1'
RG032      		ns025      		np032      		'RG2'
C032       		np032      		p          		'C2'
RG033      		ns025      		np033      		'RG3'
C033       		np033      		p          		'C3'
R030       		ns025      		ns031      		'R0'
L030       		ns031      		ns032      		'L0'
R031       		ns032      		ns033      		'R1'
L031       		ns032      		ns033      		'L1'
R032       		ns033      		ns034      		'R2'
L032       		ns033      		ns034      		'L2'
R033       		ns034      		ns035      		'R3'
L033       		ns034      		ns035      		'L3'
RG040      		ns035      		p          		'RG0'
C040       		ns035      		p          		'C0'
RG041      		ns035      		np041      		'RG1'
C041       		np041      		p          		'C1'
RG042      		ns035      		np042      		'RG2'
C042       		np042      		p          		'C2'
RG043      		ns035      		np043      		'RG3'
C043       		np043      		p          		'C3'
R040       		ns035      		ns041      		'R0'
L040       		ns041      		ns042      		'L0'
R041       		ns042      		ns043      		'R1'
L041       		ns042      		ns043      		'L1'
R042       		ns043      		ns044      		'R2'
L042       		ns043      		ns044      		'L2'
R043       		ns044      		ns045      		'R3'
L043       		ns044      		ns045      		'L3'
RG050      		ns045      		p          		'RG0'
C050       		ns045      		p          		'C0'
RG051      		ns045      		np051      		'RG1'
C051       		np051      		p          		'C1'
RG052      		ns045      		np052      		'RG2'
C052       		np052      		p          		'C2'
RG053      		ns045      		np053      		'RG3'
C053       		np053      		p          		'C3'
R050       		ns045      		ns051      		'R0'
L050       		ns051      		ns052      		'L0'
R051       		ns052      		ns053      		'R1'
L051       		ns052      		ns053      		'L1'
R052       		ns053      		ns054      		'R2'
L052       		ns053      		ns054      		'L2'
R053       		ns054      		ns055      		'R3'
L053       		ns054      		ns055      		'L3'
RG060      		ns055      		p          		'RG0'
C060       		ns055      		p          		'C0'
RG061      		ns055      		np061      		'RG1'
C061       		np061      		p          		'C1'
RG062      		ns055      		np062      		'RG2'
C062       		np062      		p          		'C2'
RG063      		ns055      		np063      		'RG3'
C063       		np063      		p          		'C3'
R060       		ns055      		ns061      		'R0'
L060       		ns061      		ns062      		'L0'
R061       		ns062      		ns063      		'R1'
L061       		ns062      		ns063      		'L1'
R062       		ns063      		ns064      		'R2'
L062       		ns063      		ns064      		'L2'
R063       		ns064      		ns065      		'R3'
L063       		ns064      		ns065      		'L3'
RG070      		ns065      		p          		'RG0'
C070       		ns065      		p          		'C0'
RG071      		ns065      		np071      		'RG1'
C071       		np071      		p          		'C1'
RG072      		ns065      		np072      		'RG2'
C072       		np072      		p          		'C2'
RG073      		ns065      		np073      		'RG3'
C073       		np073      		p          		'C3'
R070       		ns065      		ns071      		'R0'
L070       		ns071      		ns072      		'L0'
R071       		ns072      		ns073      		'R1'
L071       		ns072      		ns073      		'L1'
R072       		ns073      		ns074      		'R2'
L072       		ns073      		ns074      		'L2'
R073       		ns074      		ns075      		'R3'
L073       		ns074      		ns075      		'L3'
RG080      		ns075      		p          		'RG0'
C080       		ns075      		p          		'C0'
RG081      		ns075      		np081      		'RG1'
C081       		np081      		p          		'C1'
RG082      		ns075      		np082      		'RG2'
C082       		np082      		p          		'C2'
RG083      		ns075      		np083      		'RG3'
C083       		np083      		p          		'C3'
R080       		ns075      		ns081      		'R0'
L080       		ns081      		ns082      		'L0'
R081       		ns082      		ns083      		'R1'
L081       		ns082      		ns083      		'L1'
R082       		ns083      		ns084      		'R2'
L082       		ns083      		ns084      		'L2'
R083       		ns084      		ns085      		'R3'
L083       		ns084      		ns085      		'L3'
RG090      		ns085      		p          		'RG0'
C090       		ns085      		p          		'C0'
RG091      		ns085      		np091      		'RG1'
C091       		np091      		p          		'C1'
RG092      		ns085      		np092      		'RG2'
C092       		np092      		p          		'C2'
RG093      		ns085      		np093      		'RG3'
C093       		np093      		p          		'C3'
R090       		ns085      		ns091      		'R0'
L090       		ns091      		ns092      		'L0'
R091       		ns092      		ns093      		'R1'
L091       		ns092      		ns093      		'L1'
R092       		ns093      		ns094      		'R2'
L092       		ns093      		ns094      		'L2'
R093       		ns094      		ns095      		'R3'
L093       		ns094      		ns095      		'L3'
RG100      		ns095      		p          		'RG0'
C100       		ns095      		p          		'C0'
RG101      		ns095      		np101      		'RG1'
C101       		np101      		p          		'C1'
RG102      		ns095      		np102      		'RG2'
C102       		np102      		p          		'C2'
RG103      		ns095      		np103      		'RG3'
C103       		np103      		p          		'C3'
R100       		ns095      		ns101      		'R0'
L100       		ns101      		ns102      		'L0'
R101       		ns102      		ns103      		'R1'
L101       		ns102      		ns103      		'L1'
R102       		ns103      		ns104      		'R2'
L102       		ns103      		ns104      		'L2'
R103       		ns104      		b          		'R3'
L103       		ns104      		b          		'L3'
RG110      		b          		p          		'2*RG0'
C110       		b          		p          		'0.5*C0'
RG111      		b          		np111      		'2*RG1'
C111       		np111      		p          		'0.5*C1'
RG112      		b          		np112      		'2*RG2'
C112       		np112      		p          		'0.5*C2'
RG113      		b          		np113      		'2*RG3'
C113       		np113      		p          		'0.5*C3'
*
.ends cpw